../v/bp_fe_ras.v